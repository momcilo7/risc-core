library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package array_pkg is
	type array32 is array(natural range <>) of std_logic_vector(31 downto 0);
  	type array8 is array(natural range <>) of std_logic_vector(7 downto 0);
end package array_pkg;

package body array_pkg is
end package body array_pkg;

